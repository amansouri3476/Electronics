****************
.subckt	LPF2	1	2	0
**********input |
*****************output |
****************************GND |
L1 1 2 0.0002813
C2 2 0 5.627E-08
R3 2 0 50
.ends
