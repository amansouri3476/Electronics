****************
.subckt	LPF1	1	2	0
**********input |
*****************output |
****************************GND |
L1 1 2 0.0003751
C2 2 0 7.503E-08
R3 2 0 50
.ends
