*******************************
.subckt filter1	1	3	0
**********input |
*****************output |
****************************GND |
C1 1 2 2.001E-9
L2 2 3 562.7E-6
L1 3 0 10.00E-06
C2 3 0 112.5E-09
R8 3 0 50
.ends
