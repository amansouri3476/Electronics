****************
.subckt	HPF2	1	2	0
**********input |
*****************output |
****************************GND |
C1 1 2 225.1E-09
L2 2 0 1.125E-03
R3 2 0 50
.ends	