****************************
.subckt buffer[1]	100	200	1	4
*********************Vcc |
*****************************Vee |
**********************************input |
*****************************************output |
*************transistors
q1	100	2	3	mynpn
q2	100	3	4	mynpn
*************capacitors
c1	1	2	10u
*c2	4	5	10u
*************resistors
r1	100	2	6900k
r2	4	200	0.69k
*************models
.model	mynpn	npn	is=2f	bf=100	va=100
**************
.ends