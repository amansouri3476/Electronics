*******************************
.subckt filter2	1	3	0
**********input |
*****************output |
****************************GND |
C1 1 2 250.1E-12
L2 2 3 281.3E-6
L1 3 0 1.250E-06
C2 3 0 56.27E-09
R8 3 0 50
.ends
