****************
.subckt	HPF1	1	2	0
**********input |
*****************output |
****************************GND |
C1 1 2 1.125E-06
L2 2 0 0.005627
R3 2 0 50
.ends	