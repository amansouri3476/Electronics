****************************
.SUBCKT channel 1 2
**********input |
***********output |
E1	2	0	1	0	0.001
.ends


